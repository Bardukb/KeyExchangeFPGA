
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:13:21 12/19/2015 
// Design Name: 
// Module Name:    seg 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
module keyboarddecoder( a, seg , dig);

//input [7:0]  a;
input [3:0]  a;

output reg [6:0]dig;

output reg [3:0]seg;

always@ ( a)

begin
		seg = 4'b0000;
		case (a)
//		8'b01000101: dig <= 7'b000_0001;  // 0
//		8'b00010110: dig <= 7'b100_1111;  // 1
//		8'b00011110: dig <= 7'b001_0010;  // 2
//		8'b00100110: dig <= 7'b000_0110;  // 3
//		8'b00100101: dig <= 7'b100_1100;  // 4
//		8'b00101110: dig <= 7'b010_0100;  // 5
//		8'b00110110: dig <= 7'b010_0000;  // 6
//		8'b00111101: dig <= 7'b000_1111;  // 7
//		8'b00111110: dig <= 7'b000_0000;  // 8
//		8'b01000110: dig <= 7'b000_1100;  // 9
//		8'b00011100: dig <= 7'b000_1000;  // A
//		8'b00110010: dig <= 7'b110_0000;  // b
//		8'b00100001: dig <= 7'b111_0010;  // c
//		8'b00100011: dig <= 7'b100_0010;  // d
//		8'b00100100: dig <= 7'b011_0000;  // E
//		8'b00101011: dig <= 7'b011_1000;  // F

		4'b0000: dig <= 7'b000_0001;  // 0
		4'b0001: dig <= 7'b100_1111;  // 1
		4'b0010: dig <= 7'b001_0010;  // 2
		4'b0011: dig <= 7'b000_0110;  // 3
		4'b0100: dig <= 7'b100_1100;  // 4
		4'b0101: dig <= 7'b010_0100;  // 5
		4'b0110: dig <= 7'b010_0000;  // 6
		4'b0111: dig <= 7'b000_1111;  // 7
		4'b1000: dig <= 7'b000_0000;  // 8
		4'b1001: dig <= 7'b000_1100;  // 9
		4'b1010: dig <= 7'b000_1000;  // A
		4'b1011: dig <= 7'b110_0000;  // b
		4'b1100: dig <= 7'b111_0010;  // c
		4'b1101: dig <= 7'b100_0010;  // d
		4'b1110: dig <= 7'b011_0000;  // E
		4'b1111: dig <= 7'b011_1000;  // F

		default: dig <= 7'b111_1111 ;
		endcase		

end



endmodule

